      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "10000000100000000"; -- 1
        when "0010" => iD0 <= "10000010000010000"; -- 2
        when "0011" => iD0 <= "10001000100010000"; -- 3
        when "0100" => iD0 <= "10010001001000100"; -- 4
        when "0101" => iD0 <= "10010010010010010"; -- 5
        when "0110" => iD0 <= "10010100100101010"; -- 6
        when "0111" => iD0 <= "01010101010101010"; -- 7
        when "1000" => iD0 <= "10101010101010101"; -- 8
        when "1001" => iD0 <= "01101011011010101"; -- 9
        when "1010" => iD0 <= "01101110101101101"; -- 10
        when "1011" => iD0 <= "01101110110111011"; -- 11
        when "1100" => iD0 <= "01110111011101111"; -- 12
        when "1101" => iD0 <= "01111101111101111"; -- 13
        when "1110" => iD0 <= "01111111011111111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00000001000000001"; -- 1
        when "0010" => iD0 <= "00000100000100001"; -- 2
        when "0011" => iD0 <= "00010001000100001"; -- 3
        when "0100" => iD0 <= "00100010010001001"; -- 4
        when "0101" => iD0 <= "00100100100100101"; -- 5
        when "0110" => iD0 <= "00101001001010101"; -- 6
        when "0111" => iD0 <= "10101010101010100"; -- 7
        when "1000" => iD0 <= "01010101010101011"; -- 8
        when "1001" => iD0 <= "11010110110101010"; -- 9
        when "1010" => iD0 <= "11011101011011010"; -- 10
        when "1011" => iD0 <= "11011101101110110"; -- 11
        when "1100" => iD0 <= "11101110111011110"; -- 12
        when "1101" => iD0 <= "11111011111011110"; -- 13
        when "1110" => iD0 <= "11111110111111110"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00000010000000010"; -- 1
        when "0010" => iD0 <= "00001000001000010"; -- 2
        when "0011" => iD0 <= "00100010001000010"; -- 3
        when "0100" => iD0 <= "01000100100010010"; -- 4
        when "0101" => iD0 <= "01001001001001010"; -- 5
        when "0110" => iD0 <= "01010010010101010"; -- 6
        when "0111" => iD0 <= "01010101010101001"; -- 7
        when "1000" => iD0 <= "10101010101010110"; -- 8
        when "1001" => iD0 <= "10101101101010101"; -- 9
        when "1010" => iD0 <= "10111010110110101"; -- 10
        when "1011" => iD0 <= "10111011011101101"; -- 11
        when "1100" => iD0 <= "11011101110111101"; -- 12
        when "1101" => iD0 <= "11110111110111101"; -- 13
        when "1110" => iD0 <= "11111101111111101"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00000100000000100"; -- 1
        when "0010" => iD0 <= "00010000010000100"; -- 2
        when "0011" => iD0 <= "01000100010000100"; -- 3
        when "0100" => iD0 <= "10001001000100100"; -- 4
        when "0101" => iD0 <= "10010010010010100"; -- 5
        when "0110" => iD0 <= "10100100101010100"; -- 6
        when "0111" => iD0 <= "10101010101010010"; -- 7
        when "1000" => iD0 <= "01010101010101101"; -- 8
        when "1001" => iD0 <= "01011011010101011"; -- 9
        when "1010" => iD0 <= "01110101101101011"; -- 10
        when "1011" => iD0 <= "01110110111011011"; -- 11
        when "1100" => iD0 <= "10111011101111011"; -- 12
        when "1101" => iD0 <= "11101111101111011"; -- 13
        when "1110" => iD0 <= "11111011111111011"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00001000000001000"; -- 1
        when "0010" => iD0 <= "00100000100001000"; -- 2
        when "0011" => iD0 <= "10001000100001000"; -- 3
        when "0100" => iD0 <= "00010010001001001"; -- 4
        when "0101" => iD0 <= "00100100100101001"; -- 5
        when "0110" => iD0 <= "01001001010101001"; -- 6
        when "0111" => iD0 <= "01010101010100101"; -- 7
        when "1000" => iD0 <= "10101010101011010"; -- 8
        when "1001" => iD0 <= "10110110101010110"; -- 9
        when "1010" => iD0 <= "11101011011010110"; -- 10
        when "1011" => iD0 <= "11101101110110110"; -- 11
        when "1100" => iD0 <= "01110111011110111"; -- 12
        when "1101" => iD0 <= "11011111011110111"; -- 13
        when "1110" => iD0 <= "11110111111110111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00010000000010000"; -- 1
        when "0010" => iD0 <= "01000001000010000"; -- 2
        when "0011" => iD0 <= "00010001000010001"; -- 3
        when "0100" => iD0 <= "00100100010010010"; -- 4
        when "0101" => iD0 <= "01001001001010010"; -- 5
        when "0110" => iD0 <= "10010010101010010"; -- 6
        when "0111" => iD0 <= "10101010101001010"; -- 7
        when "1000" => iD0 <= "01010101010110101"; -- 8
        when "1001" => iD0 <= "01101101010101101"; -- 9
        when "1010" => iD0 <= "11010110110101101"; -- 10
        when "1011" => iD0 <= "11011011101101101"; -- 11
        when "1100" => iD0 <= "11101110111101110"; -- 12
        when "1101" => iD0 <= "10111110111101111"; -- 13
        when "1110" => iD0 <= "11101111111101111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00100000000100000"; -- 1
        when "0010" => iD0 <= "10000010000100000"; -- 2
        when "0011" => iD0 <= "00100010000100010"; -- 3
        when "0100" => iD0 <= "01001000100100100"; -- 4
        when "0101" => iD0 <= "10010010010100100"; -- 5
        when "0110" => iD0 <= "00100101010100101"; -- 6
        when "0111" => iD0 <= "01010101010010101"; -- 7
        when "1000" => iD0 <= "10101010101101010"; -- 8
        when "1001" => iD0 <= "11011010101011010"; -- 9
        when "1010" => iD0 <= "10101101101011011"; -- 10
        when "1011" => iD0 <= "10110111011011011"; -- 11
        when "1100" => iD0 <= "11011101111011101"; -- 12
        when "1101" => iD0 <= "01111101111011111"; -- 13
        when "1110" => iD0 <= "11011111111011111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "01000000001000000"; -- 1
        when "0010" => iD0 <= "00000100001000001"; -- 2
        when "0011" => iD0 <= "01000100001000100"; -- 3
        when "0100" => iD0 <= "10010001001001000"; -- 4
        when "0101" => iD0 <= "00100100101001001"; -- 5
        when "0110" => iD0 <= "01001010101001010"; -- 6
        when "0111" => iD0 <= "10101010100101010"; -- 7
        when "1000" => iD0 <= "01010101011010101"; -- 8
        when "1001" => iD0 <= "10110101010110101"; -- 9
        when "1010" => iD0 <= "01011011010110111"; -- 10
        when "1011" => iD0 <= "01101110110110111"; -- 11
        when "1100" => iD0 <= "10111011110111011"; -- 12
        when "1101" => iD0 <= "11111011110111110"; -- 13
        when "1110" => iD0 <= "10111111110111111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "10000000010000000"; -- 1
        when "0010" => iD0 <= "00001000010000010"; -- 2
        when "0011" => iD0 <= "10001000010001000"; -- 3
        when "0100" => iD0 <= "00100010010010001"; -- 4
        when "0101" => iD0 <= "01001001010010010"; -- 5
        when "0110" => iD0 <= "10010101010010100"; -- 6
        when "0111" => iD0 <= "01010101001010101"; -- 7
        when "1000" => iD0 <= "10101010110101010"; -- 8
        when "1001" => iD0 <= "01101010101101011"; -- 9
        when "1010" => iD0 <= "10110110101101110"; -- 10
        when "1011" => iD0 <= "11011101101101110"; -- 11
        when "1100" => iD0 <= "01110111101110111"; -- 12
        when "1101" => iD0 <= "11110111101111101"; -- 13
        when "1110" => iD0 <= "01111111101111111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00000000100000001"; -- 1
        when "0010" => iD0 <= "00010000100000100"; -- 2
        when "0011" => iD0 <= "00010000100010001"; -- 3
        when "0100" => iD0 <= "01000100100100010"; -- 4
        when "0101" => iD0 <= "10010010100100100"; -- 5
        when "0110" => iD0 <= "00101010100101001"; -- 6
        when "0111" => iD0 <= "10101010010101010"; -- 7
        when "1000" => iD0 <= "01010101101010101"; -- 8
        when "1001" => iD0 <= "11010101011010110"; -- 9
        when "1010" => iD0 <= "01101101011011101"; -- 10
        when "1011" => iD0 <= "10111011011011101"; -- 11
        when "1100" => iD0 <= "11101111011101110"; -- 12
        when "1101" => iD0 <= "11101111011111011"; -- 13
        when "1110" => iD0 <= "11111111011111110"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00000001000000010"; -- 1
        when "0010" => iD0 <= "00100001000001000"; -- 2
        when "0011" => iD0 <= "00100001000100010"; -- 3
        when "0100" => iD0 <= "10001001001000100"; -- 4
        when "0101" => iD0 <= "00100101001001001"; -- 5
        when "0110" => iD0 <= "01010101001010010"; -- 6
        when "0111" => iD0 <= "01010100101010101"; -- 7
        when "1000" => iD0 <= "10101011010101010"; -- 8
        when "1001" => iD0 <= "10101010110101101"; -- 9
        when "1010" => iD0 <= "11011010110111010"; -- 10
        when "1011" => iD0 <= "01110110110111011"; -- 11
        when "1100" => iD0 <= "11011110111011101"; -- 12
        when "1101" => iD0 <= "11011110111110111"; -- 13
        when "1110" => iD0 <= "11111110111111101"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00000010000000100"; -- 1
        when "0010" => iD0 <= "01000010000010000"; -- 2
        when "0011" => iD0 <= "01000010001000100"; -- 3
        when "0100" => iD0 <= "00010010010001001"; -- 4
        when "0101" => iD0 <= "01001010010010010"; -- 5
        when "0110" => iD0 <= "10101010010100100"; -- 6
        when "0111" => iD0 <= "10101001010101010"; -- 7
        when "1000" => iD0 <= "01010110101010101"; -- 8
        when "1001" => iD0 <= "01010101101011011"; -- 9
        when "1010" => iD0 <= "10110101101110101"; -- 10
        when "1011" => iD0 <= "11101101101110110"; -- 11
        when "1100" => iD0 <= "10111101110111011"; -- 12
        when "1101" => iD0 <= "10111101111101111"; -- 13
        when "1110" => iD0 <= "11111101111111011"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00000100000001000"; -- 1
        when "0010" => iD0 <= "10000100000100000"; -- 2
        when "0011" => iD0 <= "10000100010001000"; -- 3
        when "0100" => iD0 <= "00100100100010010"; -- 4
        when "0101" => iD0 <= "10010100100100100"; -- 5
        when "0110" => iD0 <= "01010100101001001"; -- 6
        when "0111" => iD0 <= "01010010101010101"; -- 7
        when "1000" => iD0 <= "10101101010101010"; -- 8
        when "1001" => iD0 <= "10101011010110110"; -- 9
        when "1010" => iD0 <= "01101011011101011"; -- 10
        when "1011" => iD0 <= "11011011011101101"; -- 11
        when "1100" => iD0 <= "01111011101110111"; -- 12
        when "1101" => iD0 <= "01111011111011111"; -- 13
        when "1110" => iD0 <= "11111011111110111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00001000000010000"; -- 1
        when "0010" => iD0 <= "00001000001000001"; -- 2
        when "0011" => iD0 <= "00001000100010001"; -- 3
        when "0100" => iD0 <= "01001001000100100"; -- 4
        when "0101" => iD0 <= "00101001001001001"; -- 5
        when "0110" => iD0 <= "10101001010010010"; -- 6
        when "0111" => iD0 <= "10100101010101010"; -- 7
        when "1000" => iD0 <= "01011010101010101"; -- 8
        when "1001" => iD0 <= "01010110101101101"; -- 9
        when "1010" => iD0 <= "11010110111010110"; -- 10
        when "1011" => iD0 <= "10110110111011011"; -- 11
        when "1100" => iD0 <= "11110111011101110"; -- 12
        when "1101" => iD0 <= "11110111110111110"; -- 13
        when "1110" => iD0 <= "11110111111101111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00010000000100000"; -- 1
        when "0010" => iD0 <= "00010000010000010"; -- 2
        when "0011" => iD0 <= "00010001000100010"; -- 3
        when "0100" => iD0 <= "10010010001001000"; -- 4
        when "0101" => iD0 <= "01010010010010010"; -- 5
        when "0110" => iD0 <= "01010010100100101"; -- 6
        when "0111" => iD0 <= "01001010101010101"; -- 7
        when "1000" => iD0 <= "10110101010101010"; -- 8
        when "1001" => iD0 <= "10101101011011010"; -- 9
        when "1010" => iD0 <= "10101101110101101"; -- 10
        when "1011" => iD0 <= "01101101110110111"; -- 11
        when "1100" => iD0 <= "11101110111011101"; -- 12
        when "1101" => iD0 <= "11101111101111101"; -- 13
        when "1110" => iD0 <= "11101111111011111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "00100000001000000"; -- 1
        when "0010" => iD0 <= "00100000100000100"; -- 2
        when "0011" => iD0 <= "00100010001000100"; -- 3
        when "0100" => iD0 <= "00100100010010001"; -- 4
        when "0101" => iD0 <= "10100100100100100"; -- 5
        when "0110" => iD0 <= "10100101001001010"; -- 6
        when "0111" => iD0 <= "10010101010101010"; -- 7
        when "1000" => iD0 <= "01101010101010101"; -- 8
        when "1001" => iD0 <= "01011010110110101"; -- 9
        when "1010" => iD0 <= "01011011101011011"; -- 10
        when "1011" => iD0 <= "11011011101101110"; -- 11
        when "1100" => iD0 <= "11011101110111011"; -- 12
        when "1101" => iD0 <= "11011111011111011"; -- 13
        when "1110" => iD0 <= "11011111110111111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


      case Gray0(5 downto 2) is
        when "0000" => iD0 <= "00000000000000000"; -- 0
        when "0001" => iD0 <= "01000000010000000"; -- 1
        when "0010" => iD0 <= "01000001000001000"; -- 2
        when "0011" => iD0 <= "01000100010001000"; -- 3
        when "0100" => iD0 <= "01001000100100010"; -- 4
        when "0101" => iD0 <= "01001001001001001"; -- 5
        when "0110" => iD0 <= "01001010010010101"; -- 6
        when "0111" => iD0 <= "00101010101010101"; -- 7
        when "1000" => iD0 <= "11010101010101010"; -- 8
        when "1001" => iD0 <= "10110101101101010"; -- 9
        when "1010" => iD0 <= "10110111010110110"; -- 10
        when "1011" => iD0 <= "10110111011011101"; -- 11
        when "1100" => iD0 <= "10111011101110111"; -- 12
        when "1101" => iD0 <= "10111110111110111"; -- 13
        when "1110" => iD0 <= "10111111101111111"; -- 14
        when "1111" => iD0 <= "11111111111111111"; -- 15
      end case;


